asdlfkjad